`ifndef UARTTXAGENTCONFIG_INCLUDED_
`define UARTTXAGENTCONFIG_INCLUDED_
//--------------------------------------------------------------------------------------------
// Class: UartTxAgentConfig 
// Used as the configuration class for device0 agent and it's components
//--------------------------------------------------------------------------------------------
class UartTxAgentConfig extends uvm_object;
  `uvm_object_utils(UartTxAgentConfig)

  // Variable: is_active
  // Used for creating the agent in either passive or active mode
  uvm_active_passive_enum is_active;

  //Variables
  bit hasCoverage;
  bit hasParity;
  OVER_SAMPLING_E uartOverSamplingMethod;
  BAUD_RATE_E uartBaudRate;
  DATA_TYPE_E uartDataType;/* these enum can be randomized and can apply inline constraint in test file*/
  PARITY_TYPE_E uartParityType;
  STOP_BIT_E uartStopBit;
  rand int packetsNeeded;
  bit parityErrorInjection;
//-------------------------------------------------------
// Externally defined Tasks and Functions
//-------------------------------------------------------
  extern function new(string name = "UartTxAgentConfig");

endclass : UartTxAgentConfig

//--------------------------------------------------------------------------------------------
// Construct: new
// Parameters:
// name - UartTxAgentConfig 
//--------------------------------------------------------------------------------------------
function UartTxAgentConfig :: new(string name = "UartTxAgentConfig");
  super.new(name);
endfunction : new

`endif
